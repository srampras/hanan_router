MACRO BLOCK_A
  UNITS 
    DATABASE MICRONS UNITS 1;
  END UNITS 
  ORIGIN 0 0 ;
  FOREIGN BLOCK_A 0 0 ;
  SIZE 100 BY 200 ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0 0 32 72 ;
    END
    PORT
      LAYER M3 ;
        RECT 0 0 32 72 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 64 100 96 172 ;
    END
  END B
END BLOCK_A
